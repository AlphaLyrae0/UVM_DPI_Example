`include "uvm_macros.svh"

package env_pkg;
  import uvm_pkg::*;
  import agent_pkg::*;
  import result_agent_pkg::*;
//import scoreboard_pkg::*;
//import sequence_pkg::*;
//`include "virtual_sequencer.svh"
//`include "virtual_sequence.svh"
  `include "scoreboard.svh"
  `include "env.svh"
endpackage : env_pkg
