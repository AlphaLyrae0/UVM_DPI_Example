

`include "uvm_macros.svh"

package out_agent_pkg;
  import uvm_pkg::*;
  `include "out_item.svh"
  `include "out_monitor.svh"
  `include "out_agent.svh"
endpackage
