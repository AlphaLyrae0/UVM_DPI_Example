
`include "uvm_macros.svh"

package sequence_lib_pkg;
  import uvm_pkg::*;
  import agent_pkg::*;
//import dpi_pkg::*;
//import params_pkg::*;
  `include "sequence_base.svh"
  `include "simple_sequence.svh"
  `include "dpi_sequence1.svh"
  `include "dpi_sequence2.svh"
  `include "unite_sequence.svh"
endpackage : sequence_lib_pkg
