
`include "uvm_macros.svh"

package test_lib_pkg;
  import uvm_pkg::*;
  import sequence_lib_pkg::*;
  import env_pkg::*;
  `include "test_base.svh"
  `include "simple_test.svh"
  `include "dpi_test1.svh"
  `include "dpi_test2.svh"
  `include "unite_test.svh"
endpackage : test_lib_pkg
