

`include "uvm_macros.svh"

package result_agent_pkg;
  import uvm_pkg::*;
  `include "result_item.svh"
  `include "result_monitor.svh"
  `include "result_agent.svh"
endpackage : result_agent_pkg
