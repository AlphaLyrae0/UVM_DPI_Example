
package params_pkg;
  localparam  WIDTH_p = 8;
  virtual  in_bus_if   i_vif ;
  virtual  out_bus_if  o_vif ;
endpackage : params_pkg
