`include "uvm_macros.svh"

package env_pkg;
  import uvm_pkg::*;
  import in_agent_pkg::*;
  import out_agent_pkg::*;

  `include "scoreboard.svh"
  `include "env.svh"

endpackage : env_pkg
